module cache_mem_test(cache_mem_intf.tb cmbus);

  initial
  begin : mem_t

//TO DO : Create your own stimulus (Hint call mem_write and mem_read task of cmbus instance)
  













	$finish;
  end

endmodule
